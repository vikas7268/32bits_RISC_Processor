`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.02.2020 01:01:33
// Design Name: 
// Module Name: datamem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module datamem(MemWrite,Memread,address,writeData,clk,readData);
reg[31:0] memory [0:31];
input MemWrite,Memread,clk;
input [31:0] address,writeData;
output reg [31:0] readData;
initial
begin
memory[0] = 32'b10000000000000000000000000000001;  
memory[1] = 32'b00000000000000000000000000001111;
memory[2] = 32'b00000000000000000000000000000010;
memory[3] = 32'b00000000000000000000000000000011;  
memory[4] = 32'b00000000000000000000000000000100;  
memory[5] = 32'b00000000000000000000000000000101;  
memory[6] = 32'b00000000000000000000000000000110;  
memory[7] = 32'b00000000000000000000000000000111;  
memory[8] = 32'b00000000000000000000000000001000;  
memory[9] = 32'b00000000000000000000000000001001;  
memory[10] = 32'b00000000000000000000000000001010;  
memory[11] = 32'b00000000000000000000000000001011;  
memory[12] = 32'b00000000000000000000000000001100;  
memory[13] = 32'b00000000000000000000000000001101;  
memory[14] = 32'b00000000000000000000000000000000;  
memory[15] = 32'b00000000000000000000000000000000;  
memory[16] = 32'b00000000000000000000000000000000;  
memory[17] = 32'b00000000000000000000000000000000;  
memory[18] = 32'b00000000000000000000000000000000;  
memory[19] = 32'b00000000000000000000000000000000;  
memory[20] = 32'b00000000000000000000000000000000;  
memory[21] = 32'b00000000000000000000000000000000;  
memory[22] = 32'b00000000000000000000000000000000;  
memory[23] = 32'b00000000000000000000000000000000;  
memory[24] = 32'b00000000000000000000000000000000;  
memory[25] = 32'b00000000000000000000000000000000;  
memory[26] = 32'b00000000000000000000000000000000;  
memory[27] = 32'b00000000000000000000000000000000;  
memory[28] = 32'b00000000000000000000000000000000;  
memory[29] = 32'b00000000000000000000000000000000;  
memory[30] = 32'b00000000000000000000000000000000;  
memory[31] = 32'b00000000000000000000000000000000;    
end
always@(negedge clk) 
begin
if(MemWrite==1) begin
memory[address]<=writeData;
end
end
always@(address or Memread)
begin
if(Memread==1)begin
readData=memory[address];
end
else readData=32'h0;
end
endmodule

